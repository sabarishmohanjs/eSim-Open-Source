* C:\Users\sabarishmohan\eSim-Workspace\MC14560B_test\MC14560B_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/05/25 00:06:20

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U9-Pad11_ Net-_U9-Pad12_ Net-_U9-Pad13_ Net-_U9-Pad14_ Net-_U9-Pad15_ Net-_U9-Pad16_ Net-_U10-Pad2_ Net-_U11-Pad5_ Net-_U11-Pad4_ Net-_U11-Pad3_ Net-_U11-Pad2_ Net-_U11-Pad1_ Net-_U9-Pad9_ Net-_U9-Pad10_ MC14560B		
U9  a1 b1 a2 b2 a3 b3 a4 b4 Net-_U9-Pad9_ Net-_U9-Pad10_ Net-_U9-Pad11_ Net-_U9-Pad12_ Net-_U9-Pad13_ Net-_U9-Pad14_ Net-_U9-Pad15_ Net-_U9-Pad16_ adc_bridge_8		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ adc_bridge_1		
U11  Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ Net-_U11-Pad4_ Net-_U11-Pad5_ s1 s2 s3 s4 cout dac_bridge_5		
v1  a1 GND pulse		
v3  a2 GND pulse		
v5  a3 GND pulse		
v7  a4 GND pulse		
v2  b1 GND pulse		
v4  b2 GND pulse		
v6  b3 GND pulse		
v8  b4 GND pulse		
v9  Net-_U10-Pad1_ GND DC		
U1  a1 plot_v1		
U2  b1 plot_v1		
U3  a2 plot_v1		
U4  b2 plot_v1		
U5  a3 plot_v1		
U6  b3 plot_v1		
U7  a4 plot_v1		
U8  b4 plot_v1		
U12  s1 plot_v1		
U13  s2 plot_v1		
U14  s3 plot_v1		
U15  s4 plot_v1		
U16  cout plot_v1		

.end
