* C:\Users\sabarishmohan\eSim-Workspace\54f64_test\54f64_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/22/25 14:43:48

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U2-Pad1_ Net-_U4-Pad10_ Net-_U4-Pad9_ Net-_U4-Pad8_ Net-_U4-Pad7_ Net-_U4-Pad6_ ic_54f64		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ Net-_U4-Pad5_ Net-_U4-Pad6_ Net-_U4-Pad7_ Net-_U4-Pad8_ Net-_U4-Pad9_ Net-_U4-Pad10_ adc_bridge_5		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ adc_bridge_6		
v1  Net-_U1-Pad1_ GND DC		
v2  Net-_U1-Pad2_ GND DC		
v3  Net-_U1-Pad3_ GND DC		
v4  Net-_U1-Pad4_ GND DC		
v5  Net-_U1-Pad5_ GND DC		
v6  Net-_U1-Pad6_ GND DC		
v7  Net-_U4-Pad5_ GND DC		
v8  Net-_U4-Pad4_ GND DC		
v9  Net-_U4-Pad3_ GND DC		
v10  Net-_U4-Pad2_ GND DC		
v11  Net-_U4-Pad1_ GND DC		
U2  Net-_U2-Pad1_ out dac_bridge_1		
R1  out GND 1k		
U3  out plot_v1		

.end
